library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;

entity renamer is
	port(
		a: in std_logic
	);
	
end renamer;